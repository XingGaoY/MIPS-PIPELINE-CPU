library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package cpu_pk is
type aluctr is (CT_PC,CT_LI,ct_add,ct_sub,ct_eqz,ct_eq,ct_mf,ct_nt,ct_sll,ct_srl,ct_sra,ct_or,ct_and,ct_slt,ct_un);
component alu
port(
	ctr : in aluctr;
	in1 : in std_logic_vector(15 downto 0);
	in2 : in std_logic_vector(15 downto 0);
	
	res : out std_logic_vector(15 downto 0)
	
);
end component;
component CLK_GET is
PORT(
	DYPA : OUT STD_LOGIC;
	DYPB : OUT STD_LOGIC;

	CLK : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	
	CLK36 : OUT STD_LOGIC;
	CLK18 : OUT STD_LOGIC
);
end component;
component reg is
PORT(
	REG1AD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	REG2AD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	WRREG  : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	CLK : IN STD_LOGIC;
	REGWRITEDATA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	REGWRITEADDR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CHE : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	RG1AD : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	RG2AD : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	RD1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	RD2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END component;
component SRAM
Port ( 
	DATAIN : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
   MEMMUX : in  STD_LOGIC;
   PC : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
	ADDR : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
   CLK16 : in  STD_LOGIC;
   CLK : in  STD_LOGIC;
   MEMWRT : in  STD_LOGIC;
   
	DATAOUT : out  STD_LOGIC_VECTOR(15 DOWNTO 0);
	PCPO : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	PCP : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	STALLE : IN STD_LOGIC;
	STALLO : OUT STD_LOGIC;
	
	RAM1OE : OUT STD_LOGIC;
	RAM1EN : OUT STD_LOGIC;
	RAM1WE : OUT STD_LOGIC;
	WRN : OUT STD_LOGIC;
	RDN : OUT STD_LOGIC;
	RAM1DATA : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	RAM1ADDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
	DATA_READY : in  STD_LOGIC;
   TBRE : in  STD_LOGIC;
   TSRE : in  STD_LOGIC;
	DYP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	RST : IN STD_LOGIC;
	INSTPRE : IN STD_LOGIC
);
end component;
COMPONENT IFE is
    Port ( PCP : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  PC : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
			  PCJ : in STD_LOGIC_VECTOR(15 DOWNTO 0);
           PCDT : in  STD_LOGIC;
			  PCST : IN STD_LOGIC;
           PC1 : out  STD_LOGIC_VECTOR(15 DOWNTO 0);--PC BACK TO NEXT STAGE
           PCT : out  STD_LOGIC_VECTOR(15 DOWNTO 0);--PC FOR INSTR
			  CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
			  MEM : IN STD_LOGIC;
			  IFTS : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			  DCST : OUT STD_LOGIC;
			  INSTPRE : IN STD_LOGIC);
end COMPONENT;
COMPONENT DC is
    Port ( INST : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
			  DCST : IN STD_LOGIC;
		     PCIN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);--PRESERVE THE PC FOR JUMP INSTR
			  
		     PCOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
           RD1 : out  STD_LOGIC_VECTOR(3 DOWNTO 0);
           RD2 : out  STD_LOGIC_VECTOR(3 DOWNTO 0);
           IMM : out  STD_LOGIC_VECTOR(15 DOWNTO 0);
           REGWRITE : out  STD_LOGIC;
           MEMTOREGD : out  STD_LOGIC;
           MEMWRITED : out  STD_LOGIC;
           ALUSRCD : out  STD_LOGIC;
		   
		     ALUOP_DC : OUT ALUCTR;
			  PCZERO : OUT STD_LOGIC;
			  PCJ : OUT STD_LOGIC;
		     PCOP : OUT STD_LOGIC;
		     WTREG : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		     VTMEM : OUT STD_LOGIC;
			  LWD : OUT STD_LOGIC;
			  PCST : OUT STD_LOGIC;
			  
			  STALLM : IN STD_LOGIC;
			  STALLIN : IN STD_LOGIC;
			  STALLOUT : OUT STD_LOGIC;
			  LWSTALL : IN STD_LOGIC;
			  WTREGL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  SW : OUT STD_LOGIC;
			  
			  CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
			  NUMO : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			  INSTPRE : IN STD_LOGIC;
			  INSTPREO : OUT STD_LOGIC;
			  INSTP : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  INSTPO : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		   );
end COMPONENT;
COMPONENT EXE is
    Port ( 
			  CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
			--SIGNALS FOR ALU AND PCADD
			  ALUOP : in  ALUCTR;
			  ALUSRC : in  STD_LOGIC;
			  RD1E : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  RD2E : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  IMME : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  PC : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  PCEOP : IN STD_LOGIC;
			  PCJ : IN STD_LOGIC;
			--
			--FORWARD UNIT
			  REGM : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  REGW : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  RSE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  RTE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  WREGM : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  WREGW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  RGWRITE_DE : IN STD_LOGIC;
			  REGWRITE_M : IN STD_LOGIC;
			  REGWRITE_W : IN STD_LOGIC;
			  WTREG : IN STD_LOGIC_VECTOR(3 DOWNTO 0);--
			  PCZERO_E : IN STD_LOGIC;	--	--TO CHECK IF GOTO BRANCH
			  VTMEME : IN STD_LOGIC;--
			  MEMTOREG_DE : IN STD_LOGIC;
			  MEMWRITE_DE : IN STD_LOGIC;--
			  VTMEMM : OUT STD_LOGIC;--
			  PCMUX : OUT STD_LOGIC;--
			  MEMTOREG_EM : OUT STD_LOGIC;--
			  PCE : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);--
			  RGWRITE_EM : OUT STD_LOGIC;--
			  WTREG_EM : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);--
			  ALUANS_EM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);--
			  MEMWRITE_EM : OUT STD_LOGIC;
			  RDDATA_EM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			  SW : IN STD_LOGIC;
			  SRC:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
			  );
end COMPONENT;
COMPONENT MEM is
Port ( 
	--VISIT MEM
	DATAMEM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ADDRMEM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	MEMMUX : OUT STD_LOGIC;
	MEMWRITEM : in  STD_LOGIC;
	WTMEM : OUT STD_LOGIC;	--DETERMINE TO WRITE(1) OR NOT(0)
	VTMEM : IN STD_LOGIC;	--DETERMINE WHETHER VISIT SRAM
	--
	RGWRITE_EM : in  STD_LOGIC;
   RGWRITE_MW : out  STD_LOGIC;
	RGWRITE : OUT STD_LOGIC;--DATA FOR FWU
	ALUANS_EM : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
	ALUANS_MW : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ALUANS_FWU : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
   WTREG_EM : in  STD_LOGIC_VECTOR(3 DOWNTO 0);
   WTREG_MW : out  STD_LOGIC_VECTOR(3 DOWNTO 0);
	WTREGOUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);--DATA FOR FWU
	MEMTOREG_MW : OUT STD_LOGIC;
	MEMTOREG_EM : IN STD_LOGIC;
   CLK : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	RDDATA_EM : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	MEMT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
end COMPONENT;
COMPONENT WB
	Port (
	CLK : in  STD_LOGIC;
	RST : IN STD_LOGIC;
	--DETERMINE THE DATA TO WRITE BACK
   RDMEM : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
	ALUANS_FWU : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
   ALUANS_MW : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
   DATA_W : out  STD_LOGIC_VECTOR(15 DOWNTO 0);
   MEMTOREG_MW : in  STD_LOGIC;           
	--USE TO DETERMINE FORWARD UNIT
	RGWRITE_MW : in  STD_LOGIC;
	RGWRITE_W : OUT STD_LOGIC;
   WTREG_W : out  STD_LOGIC_VECTOR(3 DOWNTO 0);
   WTREG_MW : in  STD_LOGIC_VECTOR(3 DOWNTO 0);
	WBTS : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
end COMPONENT;
end cpu_pk;