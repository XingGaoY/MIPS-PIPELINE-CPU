library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
library work;
use work.cpu_pk.all;

ENTITY REG IS
PORT(
	REG1AD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	REG2AD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	WRREG  : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	CLK : IN STD_LOGIC;
	REGWRITEDATA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	REGWRITEADDR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CHE : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	
	RG1AD : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	RG2AD : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	RD1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	RD2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	
);
END REG;

architecture reg of reg is
	TYPE RGSAVE IS ARRAY(14 DOWNTO 0) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL RG : RGSAVE;
begin
	--CHE<=WRREG&REGWRITEDATA(14 DOWNTO 0);
	CHE<=RG(8);
	PROCESS(CLK,RST)
	BEGIN
   IF(RST='0')THEN
		FOR i IN RGSAVE'RANGE LOOP
			RG(i)<=X"0000";
		END LOOP;
	ELSIF(CLK'EVENT AND CLK='0')THEN
		IF(WRREG='1')THEN
			RG(CONV_INTEGER(REGWRITEADDR))<=REGWRITEDATA;
		END IF;
	END IF;
	END PROCESS;
	
	PROCESS(CLK,REG1AD,REG2AD,RG)
	BEGIN
	IF(CLK'EVENT AND CLK='1')THEN
	IF(REG1AD/="1111")THEN
		RD1<=RG(CONV_INTEGER(REG1AD));
	ELSE
		RD1<=X"0000";
	END IF;
	IF(REG2AD/="1111")THEN
		RD2<=RG(CONV_INTEGER(REG2AD));
	ELSE
		RD2<=X"0000";
	END IF;
	RG1AD<=REG1AD;RG2AD<=REG2AD;
	END IF;
	END PROCESS;
end reg;