
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library WORK;
use WORK.CPU_PK.ALL;

entity CPU is
PORT(
	DYPA : OUT STD_LOGIC;
	DYPB : OUT STD_LOGIC;
	CLK : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	RAM1OE : OUT STD_LOGIC;
	RAM1EN : OUT STD_LOGIC;
	RAM1WE : OUT STD_LOGIC;
	WRN : OUT STD_LOGIC;
	RDN : OUT STD_LOGIC;
	RAM1DATA : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	RAM1ADDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
	DATA_READY : in  STD_LOGIC;
   TBRE : in  STD_LOGIC;
   TSRE : in  STD_LOGIC;
	LW : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	DYP1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
);
end CPU;

architecture Behavioral of CPU is
signal clk1,clk2 : std_logic;
SIGNAL PC_JUMP,PC : STD_LOGIC_VECTOR(15 DOWNTO 0);--PC VALUE FOR JUMP;
SIGNAL PC_DT : STD_LOGIC;--VALUE TO DETERMINE PC
SIGNAL PC_INS,PCIE : STD_LOGIC_VECTOR(15 DOWNTO 0);--PC FOR INSTRUCTION GET
SIGNAL LWT : STD_LOGIC;
--
SIGNAL PC_CAL : STD_LOGIC_VECTOR(15 DOWNTO 0);--PC FOR EXE STAGE TO CALCULATE NEW PC
SIGNAL PCZERO_DE,PCST : STD_LOGIC;
SIGNAL PCJ_DE : STD_LOGIC;
SIGNAL RD1_ADDR,RD2_ADDR,RSE,RTE : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL IMM_DE : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL STALL : STD_LOGIC; --STALL FOR JUMP INSTR
SIGNAL REGWRITE_DE,RGWRITE_EM,RGWRITE_MW : STD_LOGIC;
SIGNAL MEMTOREG_DE,MEMTOREG_EM,MEMTOREG_MW : STD_LOGIC;
SIGNAL MEMWRITE_DE,MEMWRITE_EM : STD_LOGIC;
SIGNAL RDDATA_EM: STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL ALUSRC_DE : STD_LOGIC;
SIGNAL ALUOP_DE : ALUCTR;
SIGNAL PCOP_DE : STD_LOGIC;
SIGNAL WTREG_DE,WTREG_EM,WTREG_MW,WTREG : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL VTMEM_DE,VTMEM_EM : STD_LOGIC;
SIGNAL REGVAL_M,REGVAL_W : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL RGDEST_M : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL RGWRITE_M,RGWRITE_W : STD_LOGIC;
SIGNAL ALUANS_EM,ALUANS_MW : STD_LOGIC_VECTOR(15 DOWNTO 0);

--
SIGNAL DATAMEM, ADDRMEM : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MEMMUX, WTMEM, SW, INSTPRE : STD_LOGIC;
SIGNAL RDMEM : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL RD1VAL, RD2VAL,INSTP : STD_LOGIC_VECTOR(15 DOWNTO 0);

SIGNAL DATA_WB : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL CHE,SRC,NUMO,IFTS,WBTS,MEMT : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL STALL1,STALL2,DCST : STD_LOGIC;
begin
LW<=SRC;
U0_clk : clk_get port map(
	DYPA => DYPA,
	DYPB => DYPB,
	CLK => clk,
	RST => rst,
	CLK36 => clk2,
	CLK18 => clk1
);
U1_IF : IFE PORT MAP(
	PCP => PC_CAL,
	PCST => PCST,
	PC => PC,
	PCJ => PC_JUMP,
   PCDT => PC_DT,
   PC1 => PC,--PC BACK TO NEXT STAGE
   PCT => PC_INS,--PC FOR INSTR
	CLK => clk2,
	RST => rst,
	MEM => MEMMUX,
	IFTS => IFTS,
	DCST => DCST,
	INSTPRE => INSTPRE
);
U2_DC : DC PORT MAP(
	INST => RDMEM,
	INSTP => INSTP,
	INSTPO => INSTP,
	DCST => DCST,
	PCIN => PCIE,--PRESERVE THE PC FOR JUMP INSTR
	PCOUT => PC_CAL,
   RD1 => RD1_ADDR,
   RD2 => RD2_ADDR,
   IMM => IMM_DE,
   REGWRITE => REGWRITE_DE,
   MEMTOREGD => MEMTOREG_DE,
   MEMWRITED => MEMWRITE_DE,
   ALUSRCD => ALUSRC_DE,
	ALUOP_DC => ALUOP_DE,
	PCOP => PCOP_DE,
	PCZERO => PCZERO_DE,
	PCJ => PCJ_DE,
	WTREG => WTREG_DE,
	VTMEM => VTMEM_DE,
	STALLM => STALL2,
	STALLIN => STALL1,
	STALLOUT => STALL1,
	LWD => LWT,
	PCST => PCST,
	LWSTALL => LWT,
	WTREGL => WTREG_DE,
	CLK => CLK2,
	RST => RST,
	NUMO => NUMO,
	INSTPRE => INSTPRE,
	INSTPREO => INSTPRE,
	SW => SW
);

U3_EXE : EXE PORT MAP(
	CLK => CLK2,
	RST => RST,
	ALUOP => ALUOP_DE,
	ALUSRC => ALUSRC_DE,
	RD1E => RD1VAL,
	RD2E => RD2VAL,
	IMME => IMM_DE,
	PC => PC_CAL,
	PCEOP => PCOP_DE,
	PCJ => PCJ_DE,
	REGM => REGVAL_M,
	REGW => REGVAL_W,
	RSE => RSE,
	RTE => RTE,
	WREGM => RGDEST_M,
	WREGW => WTREG,
	RGWRITE_DE => REGWRITE_DE,
	REGWRITE_M => RGWRITE_M,
	REGWRITE_W => RGWRITE_W, 
	WTREG => WTREG_DE,
	PCZERO_E => PCZERO_DE,	--	--TO CHECK IF GOTO BRANCH
	VTMEME => VTMEM_DE,--
	MEMTOREG_DE => MEMTOREG_DE,
	MEMWRITE_DE => MEMWRITE_DE,
	VTMEMM => VTMEM_EM,
	PCMUX => PC_DT,
	MEMTOREG_EM => MEMTOREG_EM,
	PCE => PC_JUMP,
	RGWRITE_EM => RGWRITE_EM,
	WTREG_EM => WTREG_EM,
	ALUANS_EM => ALUANS_EM,
	MEMWRITE_EM => MEMWRITE_EM,
	RDDATA_EM => RDDATA_EM,
	SW => SW,
	SRC=>SRC
);
U4_MEM : MEM PORT MAP(
	DATAMEM => DATAMEM,
	ADDRMEM => ADDRMEM,
	MEMMUX => MEMMUX,
	MEMWRITEM => MEMWRITE_EM,
	WTMEM => WTMEM,
	VTMEM => VTMEM_EM,
	--
	RGWRITE_EM => RGWRITE_EM,
   RGWRITE_MW => RGWRITE_MW,
	RGWRITE => RGWRITE_M,
	ALUANS_EM => ALUANS_EM,
	ALUANS_MW => ALUANS_MW,
	ALUANS_FWU => REGVAL_M,
   WTREG_EM => WTREG_EM,
   WTREG_MW => WTREG_MW,
	WTREGOUT => RGDEST_M,
	MEMTOREG_MW => MEMTOREG_MW,
	MEMTOREG_EM => MEMTOREG_EM,
   CLK => CLK2,
	RST => RST,
	RDDATA_EM => RDDATA_EM,
	MEMT => MEMT
);
U5_WB : WB PORT MAP(
	CLK => CLK2,
	RST => RST,
	RDMEM => RDMEM,
   DATA_W => DATA_WB,
   MEMTOREG_MW => MEMTOREG_MW,
	RGWRITE_MW => RGWRITE_MW,
	RGWRITE_W => RGWRITE_W,
   WTREG_W => WTREG,
	ALUANS_FWU => REGVAL_W,
   WTREG_MW => WTREG_MW,
	ALUANS_MW => ALUANS_MW,
	WBTS=>WBTS
);
U6_REG : REG PORT MAP(
	REG1AD => RD1_ADDR,
	REG2AD => RD2_ADDR,
	WRREG => RGWRITE_W,
	RST => RST,
	CLK => CLK2,
	REGWRITEDATA => DATA_WB,
	REGWRITEADDR => WTREG,
	RG1AD => RSE,
	RG2AD => RTE,
	RD1 => RD1VAL,
	RD2 => RD2VAL,
	CHE => CHE
);
U7_SRAM : SRAM PORT MAP(
	DATAIN => DATAMEM,
   MEMMUX => MEMMUX,
   PC =>PC_INS, 
	PCP => PC,
	PCPO => PCIE,
	ADDR => ADDRMEM,
   CLK16 => CLK,
   CLK => CLK2,
   MEMWRT => WTMEM,
	DATAOUT => RDMEM,
	STALLE =>STALL1,
	STALLO =>STALL2,
	RAM1OE => RAM1OE,
	RAM1EN => RAM1EN,
	RAM1WE => RAM1WE,
	WRN => WRN,
	RDN => RDN,
	RAM1DATA => RAM1DATA,
	RAM1ADDR => RAM1ADDR,
	DATA_READY => DATA_READY,
   TBRE => TBRE,
   TSRE => TSRE,
	DYP=> DYP1,
	RST=> RST,
	INSTPRE => INSTPRE
);
end Behavioral;

