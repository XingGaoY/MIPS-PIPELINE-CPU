
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library WORK;
use WORK.cpu_pk.all;

entity MEM is
    Port ( 
	--VISIT MEM
	DATAMEM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ADDRMEM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	MEMMUX : OUT STD_LOGIC;
	MEMWRITEM : in  STD_LOGIC;
	WTMEM : OUT STD_LOGIC;	--DETERMINE TO WRITE(1) OR NOT(0)
	VTMEM : IN STD_LOGIC;	--DETERMINE WHETHER VISIT SRAM
	--
	RGWRITE_EM : in  STD_LOGIC;
   RGWRITE_MW : out  STD_LOGIC;
	RGWRITE : OUT STD_LOGIC;--DATA FOR FWU
	ALUANS_EM : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
	ALUANS_FWU : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	RDDATA_EM : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
   WTREG_EM : in  STD_LOGIC_VECTOR(3 DOWNTO 0);
   WTREG_MW : out  STD_LOGIC_VECTOR(3 DOWNTO 0);
	WTREGOUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);--DATA FOR FWU
	MEMTOREG_MW : OUT STD_LOGIC;
	MEMTOREG_EM : IN STD_LOGIC;
   CLK : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	ALUANS_MW : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	MEMT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
end MEM;

architecture Behavioral of MEM is
begin
MEMT <= VTMEM&ALUANS_EM(15 DOWNTO 1);

RGWRITE<=RGWRITE_EM;
WTREGOUT<=WTREG_EM;
ALUANS_FWU <= ALUANS_EM;

MEMMUX<='1' WHEN(VTMEM='1')ELSE
		  '0';
WTMEM<=MEMWRITEM WHEN(RST='1')ELSE
		 '0';
ADDRMEM<=ALUANS_EM;
DATAMEM<=RDDATA_EM;

PROCESS(CLK,RST)
BEGIN
IF(RST='0')THEN
	WTREG_MW<="0000";
	RGWRITE_MW<='0';
	MEMTOREG_MW <= '0';
	ALUANS_MW <= X"0000";
ELSIF(CLK'EVENT AND CLK='1')THEN
	WTREG_MW<=WTREG_EM;
	RGWRITE_MW<=RGWRITE_EM;
	MEMTOREG_MW <= MEMTOREG_EM;
	ALUANS_MW <= ALUANS_EM;
END IF;
END PROCESS;

end Behavioral;

