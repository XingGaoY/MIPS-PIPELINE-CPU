library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library WORK;
use WORK.CPU_PK.ALL;

entity IFE is
    Port ( PCP : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  PC : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
			  PCJ : in STD_LOGIC_VECTOR(15 DOWNTO 0);
           PCDT : in  STD_LOGIC;
			  PCST : IN STD_LOGIC;
           PC1 : out  STD_LOGIC_VECTOR(15 DOWNTO 0);--PC BACK TO NEXT STAGE
           PCT : out  STD_LOGIC_VECTOR(15 DOWNTO 0);--PC FOR INSTR
			  CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
			  MEM : IN STD_LOGIC;
			  IFTS : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			  DCST : OUT STD_LOGIC;
			  INSTPRE : IN STD_LOGIC);
end IFE;

architecture IFE of IFE is
SIGNAL PCD,PC1D,PC2D,PCS : STD_LOGIC_VECTOR(15 DOWNTO 0);
begin
IFTS<=MEM&PC1D(14 DOWNTO 0);

PC2D<=PC WHEN(MEM='0')ELSE
		PC-X"0001";
		
PCS<= PCP WHEN (PCST ='1')ELSE
		PC2D;
PCD<=PCS WHEN (PCDT = '0')ELSE
	  PCJ;
	  
PC1D<=PCD+X"0001";

PROCESS(CLK,RST)
BEGIN
IF(RST='0')THEN
	PC1<=X"0000";
	PCT<=X"0000";
	DCST<='0';
ELSIF(CLK'EVENT AND CLK='1')THEN
IF(INSTPRE='1')THEN
	PC1<=PC1D-X"0001";
	PCT<=PCD-X"0001";
	DCST<=MEM;
ELSE
	PC1<=PC1D;
	PCT<=PCD;
	DCST<=MEM;
END IF;
END IF;
END PROCESS;

end IFE;

