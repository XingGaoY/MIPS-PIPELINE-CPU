library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

library WORK;
USE WORK.CPU_PK.ALL;
entity EXE is
    Port ( 
			  CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
			--SIGNALS FOR ALU AND PCADD
			  ALUOP : in  ALUCTR;
			  ALUSRC : in  STD_LOGIC;
			  RD1E : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  RD2E : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  IMME : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  PC : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  PCEOP : IN STD_LOGIC;
			  PCJ : IN STD_LOGIC;
			--
			--FORWARD UNIT
			  REGM : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  REGW : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  RSE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  RTE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  WREGM : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  WREGW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  RGWRITE_DE : IN STD_LOGIC;
			  REGWRITE_M : IN STD_LOGIC;
			  REGWRITE_W : IN STD_LOGIC;
			--
			  
			  WTREG : IN STD_LOGIC_VECTOR(3 DOWNTO 0);--
			  PCZERO_E : IN STD_LOGIC;	--	--TO CHECK IF GOTO BRANCH
			  VTMEME : IN STD_LOGIC;--
			  MEMTOREG_DE : IN STD_LOGIC;                                                        
			  MEMWRITE_DE : IN STD_LOGIC;--
			  VTMEMM : OUT STD_LOGIC;--
			  PCMUX : OUT STD_LOGIC;--
			  MEMTOREG_EM : OUT STD_LOGIC;--
			  PCE : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);--
			  RGWRITE_EM : OUT STD_LOGIC;--
			  WTREG_EM : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);--
			  ALUANS_EM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);--
			  MEMWRITE_EM : OUT STD_LOGIC;
			  RDDATA_EM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			  SW : IN STD_LOGIC;
			  
			  SRC : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
			  );
end EXE;

architecture EXE of EXE is
SIGNAL ALU2,SRCA,SRCB,PCET,RESALU:STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL FORWARDA,FORWARDB:STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL CMP,SL : STD_LOGIC;
SIGNAL ADD,IN2_ZE,SUB,SLLA,SRAA,SRLA,RDDATA : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL SHT : INTEGER;
begin
SRC<=RESALU;

IN2_ZE<=X"0000" WHEN(ALUOP=CT_EQZ)ELSE
		  SRCB;
CMP<='1' WHEN(SRCA/=IN2_ZE)ELSE
	  '0';
SL<='1' WHEN(SIGNED(SRCA)<SIGNED(IMME))ELSE
	 '0';
SHT<=8 WHEN(SRCB=X"0000")ELSE
	  TO_INTEGER(UNSIGNED(SRCB));
ADD<=STD_LOGIC_VECTOR(SIGNED(SRCA)+SIGNED(SRCB));
SUB<=STD_LOGIC_VECTOR(SIGNED(SRCA)-SIGNED(SRCB));
SLLA<=TO_STDLOGICVECTOR(TO_BITVECTOR(SRCA) SLL SHT);
SRAA<=TO_STDLOGICVECTOR(TO_BITVECTOR(SRCA) SRA SHT);
SRLA<=TO_STDLOGICVECTOR(TO_BITVECTOR(SRCA) SRL SHT);


RESALU<=ADD 								WHEN(ALUOP=CT_ADD)ELSE
	  SUB									WHEN(ALUOP=CT_SUB)ELSE
	  SRCA AND SRCB 						WHEN(ALUOP=CT_AND)ELSE
	  SRCA									WHEN(ALUOP=CT_MF)ELSE
	  NOT SRCA							WHEN(ALUOP=CT_NT)ELSE
	  SRCA OR SRCB						WHEN(ALUOP=CT_OR)ELSE
	  SLLA								WHEN(ALUOP=CT_SLL)ELSE
	  SRAA								WHEN(ALUOP=CT_SRA)ELSE
	  SRLA								WHEN(ALUOP=CT_SRL)ELSE
	  (0=>SL,OTHERS=>'0')			WHEN(ALUOP=CT_SLT)ELSE
	  (0=>CMP,OTHERS=>'0')			WHEN((ALUOP=CT_EQZ)OR(ALUOP=CT_EQ))ELSE
	  SRCB								WHEN(ALUOP=CT_LI)ELSE
	  PC									WHEN(ALUOP=CT_PC)ELSE
	  (OTHERS=>'0');
PROCESS(CLK,RST)
BEGIN
IF(RST='0')THEN
	MEMWRITE_EM<='0';
	VTMEMM<='0';
	RGWRITE_EM<='0';
	WTREG_EM<=X"0";
	MEMTOREG_EM<='0';
--	PCE<=X"0000";
	ALUANS_EM<=X"0000";
	RDDATA_EM<=X"0000";
ELSIF(CLK'EVENT AND CLK='1')THEN
	MEMWRITE_EM<=MEMWRITE_DE;
	VTMEMM<=VTMEME;
	RGWRITE_EM<=RGWRITE_DE;
	MEMTOREG_EM<=MEMTOREG_DE;
	WTREG_EM<=WTREG;
--	PCE<=PCET;
	ALUANS_EM<=RESALU;
	RDDATA_EM<=RDDATA;
END IF;
END PROCESS;

PCE<=STD_LOGIC_VECTOR(SIGNED(PC)+SIGNED(IMME)) WHEN(PCEOP='1')AND(RST='1') ELSE
	  RD1E WHEN(PCEOP='0')AND(RST='1')ELSE
	  X"0000";

ALU2<=RD2E WHEN(ALUSRC='0')ELSE
	   IMME;
		
RDDATA <= REGM WHEN ((RTE/="1111") AND (RTE=WREGM) AND (REGWRITE_M='1')) ELSE
			 REGW WHEN ((RTE/="1111") AND (RTE=WREGW) AND (REGWRITE_W='1')) ELSE
			 RD2E;

FORWARDA<="10" WHEN ((RSE/="1111") AND (RSE=WREGM) AND (REGWRITE_M='1')) ELSE
		    "01" WHEN ((RSE/="1111") AND (RSE=WREGW) AND (REGWRITE_W='1')) ELSE
		    "00";
		  
FORWARDB<="10" WHEN ((RTE/="1111") AND (RTE=WREGM) AND (REGWRITE_M='1')) ELSE
		    "01" WHEN ((RTE/="1111") AND (RTE=WREGW) AND (REGWRITE_W='1')) ELSE
		    "00";
		  
SRCA <= RD1E WHEN(FORWARDA="00")ELSE
	     REGW WHEN(FORWARDA="01")ELSE
	     REGM WHEN(FORWARDA="10")ELSE
	     X"0000";
	  
SRCB <= ALU2 WHEN(FORWARDB="00")OR(SW='1')ELSE
	     REGW WHEN(FORWARDB="01")AND(SW='0')ELSE
	     REGM WHEN(FORWARDB="10")AND(SW='0')ELSE
	     X"0000";
		  
PCMUX<='1'WHEN(((PCJ='1')AND(PCZERO_E='0')AND(RESALU(0)='0'))OR((PCJ='1')AND(PCZERO_E='1')AND(RESALU(0)='1')))ELSE
		 '0';

end EXE;

