library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library WORK;
use WORK.cpu_pk.all;

entity DC is
    Port ( INST : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
			  INSTP : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			  INSTPO : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			  DCST : IN STD_LOGIC;
		     PCIN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);--PRESERVE THE PC FOR JUMP INSTR
			  
		     PCOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
           RD1 : out  STD_LOGIC_VECTOR(3 DOWNTO 0);
           RD2 : out  STD_LOGIC_VECTOR(3 DOWNTO 0);
           IMM : out  STD_LOGIC_VECTOR(15 DOWNTO 0);
           REGWRITE : out  STD_LOGIC;
           MEMTOREGD : out  STD_LOGIC;
           MEMWRITED : out  STD_LOGIC;
           ALUSRCD : out  STD_LOGIC;
		   
		     ALUOP_DC : OUT ALUCTR;
			  PCZERO : OUT STD_LOGIC;
			  PCJ : OUT STD_LOGIC;
		     PCOP : OUT STD_LOGIC;
		     WTREG : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		     VTMEM : OUT STD_LOGIC;
			  LWD : OUT STD_LOGIC;
			  PCST : OUT STD_LOGIC;
			  
			  STALLIN : IN STD_LOGIC;
			  STALLM : IN STD_LOGIC;
			  STALLOUT : OUT STD_LOGIC;
			  LWSTALL : IN STD_LOGIC;
			  WTREGL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  SW : OUT STD_LOGIC;
			  
			  CLK : IN STD_LOGIC;
			  RST : IN STD_LOGIC;
			  INSTPREO : OUT STD_LOGIC;
			  INSTPRE : IN STD_LOGIC;
			  NUMO : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		   );
end DC;

architecture DC of DC is
TYPE IMMTP IS(IMM10,IMM7,IMM4,IMM3,IMMSL,IMMZE,IMMNON);
TYPE INS IS
RECORD
OP : STD_LOGIC_VECTOR(9 DOWNTO 0);
CTR : ALUCTR;
RSP : STD_LOGIC_VECTOR(2 DOWNTO 0);--"000"ONE REG,"001"TWO TEG,"010"ONE SP REG,"011"TWO REG WITH ONE SP,"100"NO REG
RREGPS : STD_LOGIC_VECTOR(3 DOWNTO 0);--IF SP_REG='0'AND REGPS=0xF CHOOSE RD2T TO BE RD1A, ELSE RD1T OR THE SPREG
WSP_REG : STD_LOGIC_VECTOR(1 DOWNTO 0);--"00"RG,"01"RSP,"10"NORG
RDESTD : STD_LOGIC_VECTOR(3 DOWNTO 0);--0x0 WHEN RD1, 0x1 WHEN RD2,Ox2 WHEN RD3,0xSP
WRITEREG : STD_LOGIC;
IMMTYPE : IMMTP;
SRC : STD_LOGIC;
PCE : STD_LOGIC;
PCZR : STD_LOGIC;
PCJ : STD_LOGIC;
MEM : STD_LOGIC;
MEMW : STD_LOGIC;
ALUSR : STD_LOGIC;
MEMTOR : STD_LOGIC;
SW : STD_LOGIC;
END RECORD;
SIGNAL INSRPS : INTEGER RANGE 0 TO 29;
SIGNAL LW,STALL,PCS,CON_ST : STD_LOGIC;
SIGNAL STALLT : STD_LOGIC;
SIGNAL RDST : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL IMMT1,INSTT : STD_LOGIC_VECTOR(15 DOWNTO 0);
TYPE INS_TYPE IS ARRAY (0 TO 29)OF INS;
CONSTANT INS_TABLE : INS_TYPE :=
(
--INSTRUCTION TABLE
("0100100000",CT_ADD,"000","0000","00","0000",'1',IMM7,'1','0','0','0','0','0','1','0','0'),--ADD
("0100000000",CT_ADD,"000","0000","00","0001",'1',IMM3,'1','0','0','0','0','0','1','0','0'),--ADDIU3
("0110001100",CT_ADD,"010","1000","01","1000",'1',IMM7,'1','0','0','0','0','0','1','0','0'),--ADDSP
("1110001000",CT_ADD,"001","0000","00","0010",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--ADDU
("1110101100",CT_AND,"001","0000","00","0000",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--AND
("0001000000",CT_UN, "100","0000","10","0000",'0',IMM10,'1','1','0','1','0','0','0','0','0'),--B
("0010000000",CT_EQZ,"000","0000","10","0000",'0',IMM7,'1','1','0','1','0','0','0','0','0'),--BEQZ
("0010100000",CT_EQZ,"000","0000","10","0000",'0',IMM7,'1','1','1','1','0','0','0','0','0'),--BNEZ
("0110000000",CT_EQZ,"010","1001","10","0000",'0',IMM7,'1','1','0','1','0','0','0','0','0'),--BTEQZ
("1110101010",CT_EQ, "001","0000","01","1001",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--CMP
("0111000000",CT_EQ, "000","0000","01","1001",'1',IMM7,'1','0','0','0','0','0','1','0','0'),--CMPI
("1110100000",CT_UN, "000","0000","10","0000",'0',IMMNON,'0','0','0','1','0','0','0','0','0'),--JR
("0110100000",CT_LI, "000","0000","00","0000",'1',IMMZE,'1','0','0','0','0','0','1','0','0'),--LI
("1001100000",CT_ADD,"000","0000","00","0001",'1',IMM4,'1','0','0','0','1','0','1','1','0'),--LW
("1001000000",CT_ADD,"010","1000","00","0000",'1',IMM7,'1','0','0','0','1','0','1','1','0'),--LW_SP
("1111000000",CT_MF, "010","1010","00","0000",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--MFIH
("1110110000",CT_PC, "100","0000","00","0000",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--MFPC
("0111100000",CT_MF, "000","1111","00","0000",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--MOVE
("1111010000",CT_MF, "000","0000","01","1010",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--MTIH
("0110010000",CT_MF, "000","1111","01","1000",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--MTSP
("1110101111",CT_NT,"000","1111","00","0000",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--NOT
("1110101101",CT_OR, "001","0000","00","0000",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--OR
("0000100000",CT_UN, "100","0000","10","0000",'0',IMMNON,'0','0','0','0','0','0','0','0','0'),--NOP
("0011000000",CT_SLL,"000","1111","00","0000",'1',IMMSL,'1','0','0','0','0','0','1','0','0'),--SLL
("0101000000",CT_SLT,"000","0000","01","1001",'1',IMM7,'1','0','0','0','0','0','1','0','0'),--SLTI
("0011011000",CT_SRA,"000","1111","00","0000",'1',IMMSL,'1','0','0','0','0','0','1','0','0'),--SRA
("0011010000",CT_SRL,"000","1111","00","0000",'1',IMMSL,'1','0','0','0','0','0','1','0','0'),--SRL
("1110011000",CT_SUB,"001","0000","00","0010",'1',IMMNON,'0','0','0','0','0','0','0','0','0'),--SUBU
("1101100000",CT_ADD,"001","0000","10","0000",'0',IMM4,'1','0','0','0','1','1','1','0','1'),--SW
("1101000000",CT_ADD,"011","1000","10","0000",'0',IMM7,'1','0','0','0','1','1','1','0','0')--SW_SP
);
begin
INSTT<=INST WHEN INSTPRE='0' ELSE
		 INSTP;
PROCESS(INSTT,LWSTALL,WTREGL)
VARIABLE IMMT:STD_LOGIC_VECTOR(15 DOWNTO 0);
VARIABLE INS_OP : STD_LOGIC_VECTOR(9 DOWNTO 0);
VARIABLE UN_INS : STD_LOGIC;
VARIABLE NUM : INTEGER RANGE 0 TO 30;
VARIABLE RD1T,RD2T,RD3T,RD1T1,RD2T1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
IF(INSTT(15 DOWNTO 11)="11101")THEN
	IF(INSTT(4 DOWNTO 0)="00000")THEN
		INS_OP := INSTT(15 DOWNTO 11)&INSTT(6 DOWNTO 2);
	ELSE
		INS_OP := INSTT(15 DOWNTO 11)&INSTT(4 DOWNTO 0);
	END IF;
ELSIF(INSTT(15 DOWNTO 11)="01100")THEN
INS_OP := INSTT(15 DOWNTO 8)&"00";
ELSIF(INSTT(15 DOWNTO 11)="11100")THEN
INS_OP := INSTT(15 DOWNTO 11)&INSTT(1 DOWNTO 0)&"000";
ELSIF(INSTT(15 DOWNTO 11)="00110")THEN
INS_OP := INSTT(15 DOWNTO 11)&INSTT(1 DOWNTO 0)&"000";
ELSIF(INSTT(15 DOWNTO 11)="11110")THEN
INS_OP := INSTT(15 DOWNTO 11)&INSTT(0)&"0000";
ELSE
INS_OP := INSTT(15 DOWNTO 11)&"00000";
END IF;
UN_INS := '0';
FOR i IN INS_TABLE'RANGE LOOP
	IF INS_TABLE(i).OP=INS_OP THEN
		UN_INS:='1';
		NUM:=i;
		EXIT;
	ELSE
		NUM:=30;
	END IF;
END LOOP;
INSRPS<=NUM;
NUMO<=CONV_STD_LOGIC_VECTOR(NUM,16);
IF(NUM=13)OR(NUM=14)THEN
LW<='1';
ELSE
LW<='0';
END IF;

RD1T:='0'&INSTT(10 DOWNTO 8);
RD2T:='0'&INSTT(7 DOWNTO 5);
RD3T:='0'&INSTT(4 DOWNTO 2);

IF((INS_TABLE(NUM).RSP="000")AND(INS_TABLE(NUM).RREGPS="0000"))THEN
	RD1T1:=RD1T;RD2T1:="1111";
ELSIF((INS_TABLE(NUM).RSP="000")AND(INS_TABLE(NUM).RREGPS="1111"))THEN
	RD1T1:=RD2T;RD2T1:="1111";
ELSIF((INS_TABLE(NUM).RSP="001"))THEN
	RD1T1:=RD1T;RD2T1:=RD2T;
ELSIF((INS_TABLE(NUM).RSP)="010")THEN
	RD1T1:=INS_TABLE(NUM).RREGPS;RD2T1:="1111";
ELSIF(INS_TABLE(NUM).RSP="011")THEN
	RD1T1:=INS_TABLE(NUM).RREGPS;RD2T1:=RD1T;
ELSE
	RD1T1:="1111";RD2T1:="1111";
END IF;
RD1<=RD1T1;RD2<=RD2T1;
IF(INS_TABLE(NUM).WSP_REG="00")THEN
	CASE INS_TABLE(NUM).RDESTD IS
	WHEN "0000"=>RDST<=RD1T;
	WHEN "0001"=>RDST<=RD2T;
	WHEN "0010"=>RDST<=RD3T;
	WHEN OTHERS=>RDST<=X"0";
	END CASE;
ELSIF(INS_TABLE(NUM).WSP_REG="01")THEN
	RDST<=INS_TABLE(NUM).RDESTD;
ELSE
	RDST<="1011";
END IF;

IF((NUM=5)OR(NUM=6)OR(NUM=7)OR(NUM=8)OR(NUM=11))THEN
STALL<='1';PCS<='1';
ELSE
STALL<='0';PCS<='0';
END IF;

IF(LWSTALL='1')AND((WTREGL=RD1T1)OR(WTREGL=RD2T1))THEN
CON_ST<='1';
ELSE
CON_ST<='0';
END IF;

CASE INS_TABLE(NUM).IMMTYPE IS
WHEN IMM10=>
	IF(INSTT(10)='0')THEN
		IMMT:="00000"&INSTT(10 DOWNTO 0);
	ELSE
		IMMT:="11111"&INSTT(10 DOWNTO 0);
	END IF;
WHEN IMM7=>
	IF(INSTT(7)='0')THEN
		IMMT:="00000000"&INSTT(7 DOWNTO 0);
	ELSE
		IMMT:="11111111"&INSTT(7 DOWNTO 0);
	END IF;
WHEN IMM4=>
	IF(INSTT(4)='0')THEN
		IMMT:="00000000000"&INSTT(4 DOWNTO 0);
	ELSE
		IMMT:="11111111111"&INSTT(4 DOWNTO 0);
	END IF;
WHEN IMM3=>
	IF(INSTT(3)='0')THEN
		IMMT:="000000000000"&INSTT(3 DOWNTO 0);
	ELSE
		IMMT:="111111111111"&INSTT(3 DOWNTO 0);
	END IF;
WHEN IMMSL=>
	IF(INSTT(4)='0')THEN
		IMMT:="0000000000000"&INSTT(4 DOWNTO 2);
	ELSE							
		IMMT:="1111111111111"&INSTT(4 DOWNTO 2);
	END IF;
WHEN IMMZE=>
	IMMT:="00000000"&INSTT(7 DOWNTO 0);
WHEN IMMNON=>
	IMMT:=X"0000";
END CASE;
IMMT1<=IMMT;
END PROCESS;

STALLT<=STALLIN OR STALLM;

PROCESS(CLK,RST)
BEGIN
IF(RST='0')THEN
	ALUOP_DC<=CT_UN;
	IMM<=X"0000";
	PCOUT<=X"0000";
	PCOP<='0';	
	REGWRITE<='0';
	WTREG<=X"0";
	VTMEM<='0';
	PCZERO <= '0';
	PCJ <= '0';
	MEMWRITED <= '0';
	STALLOUT <= '0';
	LWD<='0';
	ALUSRCD<='0';
	MEMTOREGD<='0';
	PCST<='0';
	SW<='0';
	INSTPREO<='0';
	INSTPO<=X"0000";
	
ELSIF(CLK'EVENT AND CLK='1')THEN
IF(INSTT=X"0000")OR(STALLT='1')OR(INSRPS=30)OR(DCST='1')THEN
	ALUOP_DC<=CT_UN;
	IMM<=X"0000";
	PCOUT<=X"0000";
	PCOP<='0';	
	REGWRITE<='0';
	WTREG<=X"0";
	VTMEM<='0';
	PCZERO <= '0';
	PCJ <= '0';
	MEMWRITED <= '0';
	STALLOUT <= '0';
	LWD<='0';
	ALUSRCD<='0';
	MEMTOREGD<='0';
	PCST<='0';
	SW<='0';
	INSTPREO<='0';
	INSTPO<=X"0000";
ELSIF CON_ST='1' THEN
	ALUOP_DC<=CT_UN;
	IMM<=X"0000";
	PCOUT<=X"0000";
	PCOP<='0';	
	REGWRITE<='0';
	WTREG<=X"0";
	VTMEM<='0';
	PCZERO <= '0';
	PCJ <= '0';
	MEMWRITED <= '0';
	STALLOUT <= '0';
	LWD<='0';
	ALUSRCD<='0';
	MEMTOREGD<='0';
	PCST<='0';
	SW<='0';
	INSTPREO<='1';
	INSTPO<=INST;
ELSE
	ALUOP_DC<=INS_TABLE(INSRPS).CTR;
	IMM<=IMMT1;
	PCOUT<=PCIN;
	PCOP<=INS_TABLE(INSRPS).PCE;
	REGWRITE <= INS_TABLE(INSRPS).WRITEREG;
	WTREG<=RDST;
	VTMEM<=INS_TABLE(INSRPS).MEM;
	PCZERO <= INS_TABLE(INSRPS).PCZR;
	PCJ <= INS_TABLE(INSRPS).PCJ;
	MEMWRITED <= INS_TABLE(INSRPS).MEMW;
	STALLOUT<=STALL;
	LWD<=LW;
	ALUSRCD<=INS_TABLE(INSRPS).ALUSR;
	MEMTOREGD<=INS_TABLE(INSRPS).MEMTOR;
	PCST<=PCS;
	SW<=INS_TABLE(INSRPS).SW;
	INSTPREO<='0';
	INSTPO<=X"0000";
END IF;
END IF;
END PROCESS;

end DC;

