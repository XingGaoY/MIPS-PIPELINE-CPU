library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library WORK;
USE WORK.CPU_PK.ALL;

entity WB is
    Port ( CLK : in  STD_LOGIC;
			  RST : IN STD_LOGIC;
	
		--DETERMINE THE DATA TO WRITE BACK
           RDMEM : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
           ALUANS_MW : in  STD_LOGIC_VECTOR(15 DOWNTO 0);
           DATA_W : out  STD_LOGIC_VECTOR(15 DOWNTO 0);
           MEMTOREG_MW : in  STD_LOGIC;           
		--USE TO DETERMINE FORWARD UNIT
			  RGWRITE_MW : in  STD_LOGIC;
		     RGWRITE_W : OUT STD_LOGIC;
           WTREG_W : out  STD_LOGIC_VECTOR(3 DOWNTO 0);
           WTREG_MW : in  STD_LOGIC_VECTOR(3 DOWNTO 0);
			  ALUANS_FWU : out STD_LOGIC_VECTOR(15 DOWNTO 0);
			  WBTS : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
			  );
end WB;

architecture WB of WB is	
SIGNAL DATA : STD_LOGIC_VECTOR(15 DOWNTO 0);
begin
WBTS<=DATA;
DATA<=RDMEM WHEN(MEMTOREG_MW = '1')ELSE
		ALUANS_MW;
DATA_W <= DATA;
WTREG_W<=WTREG_MW;
RGWRITE_W<=RGWRITE_MW WHEN(RST='1')ELSE
		  '0';
ALUANS_FWU <= DATA;
end WB;

